// pipelined MIPS processor
module mipspipe(input logic clk, reset,
	    output logic [31:0] pcF,
	    input logic [31:0] instrF,
 	    output logic memwriteM,
	    output logic [31:0] aluoutM, writedataM,
	    input logic [31:0] readdataM);

	logic [5:0] opD, functD;
	logic [1:0] memtoregE, memtoregM, memtoregW;
	logic regdstE, alusrcE,pcsrcD,regwriteE, regwriteM, regwriteW;
	logic [3:0] alucontrolE;
	logic flushE, equalD;
	logic sbE, sbM, lbE, lbM, lbW,jalregW;

	controllerpipe c(clk, reset, opD, functD, flushE,
			equalD,memtoregE, memtoregM,
			memtoregW, memwriteM, pcsrcD,
			branchD, bneD, alusrcE, regdstE, regwriteE,
			regwriteM, regwriteW, jumpD, jrD, jalD, jalE,jalregE, jalregM, jalregW,
			alucontrolE, sbE, sbM, lbE, lbM, lbW);

	datapathpipe dp(clk, reset, memtoregE, memtoregM,
		        memtoregW, pcsrcD, branchD, bneD,
			alusrcE, regdstE, regwriteE,
			regwriteM, regwriteW, jumpD, jrD,sbM, lbW, jalD, jalE,jalregW, 
			alucontrolE,
			equalD, pcF, instrF,
			aluoutM, writedataM, readdataM,
			opD, functD, flushE);

endmodule


module  controllerpipe (input logic clk, reset,
			input logic [5:0] opD, functD,
			input logic flushE, equalD,
			output logic [1:0] memtoregE,memtoregM, memtoregW,
			output logic memwriteM,
			output logic pcsrcD,branchD, bneD, alusrcE,
			output logic regdstE,regwriteE,
			output logic regwriteM,regwriteW,
			output logic jumpD, jrD, jalD, jalE, jalregE, jalregM, jalregW,
			output logic [3:0] alucontrolE,
			output logic sbE, sbM,lbE, lbM, lbW);

		logic [1:0] aluopD, memtoregD;
		logic  memwriteD, alusrcD,regdstD, regwriteD;
		logic [3:0] alucontrolD;
		logic memwriteE;
		logic sbD, lbD,jalregD;

	maindecpipe md(opD, functD, memtoregD, memwriteD, branchD, bneD, alusrcD, regdstD, regwriteD, jumpD, jrD, jalD, aluopD, sbD, lbD,jalregD);

	aludecpipe ad(functD, aluopD, alucontrolD);

	assign pcsrcD = (branchD & equalD) | (bneD & ~equalD);

// pipeline registers
	floprc #(14) regE(clk, reset, flushE,
			{memtoregD, memwriteD, alusrcD,regdstD, regwriteD, alucontrolD, sbD, lbD, jalD,jalregD},
			{memtoregE, memwriteE, alusrcE,regdstE, regwriteE, alucontrolE, sbE, lbE, jalE,jalregE});

	flopr #(7) regM(clk, reset,
			{memtoregE, memwriteE, regwriteE, sbE, lbE,jalregE},
			{memtoregM, memwriteM, regwriteM, sbM, lbM,jalregM});

	flopr #(5) regW(clk, reset,
			{memtoregM, regwriteM, lbM, jalregM},
			{memtoregW, regwriteW, lbW, jalregW});

endmodule


module maindecpipe(input logic [5:0] op, funct,
		output logic [1:0] memtoreg,
		output logic memwrite, branch, bne, alusrc,
		output logic regdst, regwrite,
		output logic jump, jr, jal,
		output logic [1:0] aluop,
		output logic sb, lb, jalreg);

	logic [15:0] controls;
	assign {regwrite, regdst, alusrc,branch, bne, memwrite,memtoreg, jump, aluop, sb, lb, jr, jal,jalreg} = controls;
//here
	always_comb
	case(op)
	6'b000000: 
		case(funct)
		6'b010010: controls <= 16'b1100001001000000; //mflo
		6'b010000: controls <= 16'b1100001101000000; //mfhi
		6'b001000: controls <= 16'b1100000001000100; //jr
		default:   controls <= 16'b1100000001000000; //Rtyp
		endcase

	6'b100011: controls <= 16'b1010000100000000; //LW
	6'b101011: controls <= 16'b0010010000000000; //SW
	6'b000100: controls <= 16'b0001000000100000; //BEQ
	6'b001000: controls <= 16'b1010000000000000; //ADDI
	6'b000010: controls <= 16'b0000000010000000; //J
	6'b000101: controls <= 16'b0000100000100000; //bne
	6'b001010: controls <= 16'b1010000001100000; //slti
	6'b101000: controls <= 16'b0010010000010000; //sb
	6'b100000: controls <= 16'b1010000100001000; //lb
	6'b001000: controls <= 16'b1100000001000100; //jr
	6'b000011: controls <= 16'b0000000010000011; //jal
	default: controls <= 16'bxxxxxxxxxxxxxxxx; //???
	endcase
endmodule



module aludecpipe(input logic [5:0] funct,
	input logic [1:0] aluop,
	output logic [3:0] alucontrol);
//here
	always_comb
	case(aluop)
	2'b00: alucontrol <= 4'b0010; // add
	2'b01: alucontrol <= 4'b0110; // sub
	2'b11: alucontrol <= 4'b0111; //slti
	default: case(funct) // RTYPE
		6'b100000: alucontrol <= 4'b0010; // ADD
		6'b100010: alucontrol <= 4'b0110; // SUB
		6'b100100: alucontrol <= 4'b0000; // AND
		6'b100101: alucontrol <= 4'b0001; // OR
		6'b101010: alucontrol <= 4'b0111; // SLT
		6'b011000: alucontrol <= 4'b1010; //multiply
		6'b011010: alucontrol <= 4'b1011; //division
		6'b000000: alucontrol <= 4'b1000; //shift left logical
		6'b000010: alucontrol <= 4'b1001; //shift right logical
		default: alucontrol <= 4'bxxxx; // ???
		endcase
	endcase
endmodule


module datapathpipe(input logic clk, reset,
		input logic [1:0] memtoregE,memtoregM,memtoregW,
		input logic pcsrcD, branchD, bneD,
		input logic alusrcE, regdstE,
		input logic regwriteE,regwriteM,regwriteW,
		input logic jumpD, jrD, sbM, lbW, jalD, jalE,jalregW,
		input logic [3:0] alucontrolE,
		output logic equalD,
		output logic [31:0] pcF,
		input logic [31:0] instrF,
		output logic [31:0] aluoutM,writedataM,
		input logic [31:0] readdataM,
		output logic [5:0] opD, functD,
		output logic flushE);

	logic forwardaD, forwardbD;
	logic [1:0] forwardaE, forwardbE;
	logic stallF;
	logic [4:0] rsD, rtD, rdD, rsE, rtE, rdE;
	logic [4:0] writeregE, writeregM, writeregW,temp;
	logic flushD;
	logic [31:0] pcnextFD, pcnextbrFD,pcplus4F, pcbranchD, pcplus4E, pcplus4M, pcplus4W;
	logic [31:0] signimmD, signimmE, signimmshD;
	logic [31:0] srcaD, srca2D, srcaE, srca2E;
	logic [31:0] srcbD, srcb2D, srcbE, srcb2E, srcb3E;
	logic [31:0] pcplus4D, instrD,instrE, instrM, instrW;
	logic [31:0] aluoutE, aluoutW;
	logic [31:0] readdataW, resultW;
//here
	logic [31:0] lo, hi, loM, loW, hiM, hiW,hiE,loE;
	logic [63:0] m;
	logic [4:0] shamtD, shamtE;
	logic [7:0] lbyte, sbyte;
	logic [31:0] exlbyte, exsbyte;
	

	
	
// hazard detection
	hazard h(rsD, rtD, rsE, rtE, writeregE, writeregM,writeregW,regwriteE, regwriteM, regwriteW,memtoregE, memtoregM, branchD, bneD, forwardaD, forwardbD, forwardaE,forwardbE,stallF, stallD, flushE);

// register file (operates in decode and writeback)
	regfilepipe rf(clk, regwriteW, rsD, rtD, writeregW,resultW, srcaD, srcbD);


// next PC logic (operates in fetch and decode)
	mux2 #(32) pcbrmux(pcplus4F, pcbranchD, pcsrcD,pcnextbrFD);
	mux2 #(32) pcmux(pcnextbrFD,{pcplus4D[31:28],instrD[25:0], 2'b00},jumpD, pcnextFD);
	mux2 #(32) pcjr(pcnextFD, srca2D, jrD, pcnextFD);

// Fetch stage logic
	flopenr #(32) pcreg(clk, reset, ~stallF,pcnextFD, pcF);
	adder pcadd1(pcF, 32'b100, pcplus4F);

// Decode stage
	flopenr #(32) r1D(clk, reset, ~stallD, pcplus4F,pcplus4D);
	flopenrc #(32) r2D(clk, reset, ~stallD, flushD, instrF,instrD);
	

	signext se(instrD[15:0], signimmD);
	sl2 immsh(signimmD, signimmshD);
	adder pcadd2(pcplus4D, signimmshD, pcbranchD);
	mux2 #(32) forwardadmux(srcaD, aluoutM, forwardaD,srca2D);
	mux2 #(32) forwardbdmux(srcbD, aluoutM, forwardbD,srcb2D);
	eqcmp comp(srca2D, srcb2D, equalD);

//here
	assign shamtD = instrD[10:6];
	assign opD = instrD[31:26];
	assign functD = instrD[5:0];
	assign rsD = instrD[25:21];
	assign rtD = instrD[20:16];
	assign rdD = instrD[15:11];
	assign flushD = pcsrcD | jumpD | jrD;
// Execute stage
	floprc #(32) r1E(clk, reset, flushE, srcaD, srcaE);
	floprc #(32) r2E(clk, reset, flushE, srcbD, srcbE);
	floprc #(32) r3E(clk, reset, flushE, signimmD, signimmE);
	floprc #(32) pc1(clk, reset, flushE, pcplus4D, pcplus4E);
	floprc #(32) instr1(clk, reset, flushE, instrD, instrE);
	floprc #(5) r4E(clk, reset, flushE, rsD, rsE);
	floprc #(5) r5E(clk, reset, flushE, rtD, rtE);
	floprc #(5) r6E(clk, reset, flushE, rdD, rdE);
	floprc #(5) shamt(clk, reset, flushE, shamtD, shamtE);
//here
	
	mux3 #(32) forwardaemux(srcaE, resultW, aluoutM,forwardaE, srca2E);
	mux3 #(32) forwardbemux(srcbE, resultW, aluoutM,forwardbE, srcb2E);
	mux2 #(32) srcbmux(srcb2E, signimmE, alusrcE,srcb3E);
//here
	ALUpipeall alu(srca2E, srcb3E, alucontrolE, shamtE, aluoutE, hi, lo, m);
	mux2 #(5) wrmux(rtE, rdE, regdstE, temp);
	mux2 #(5) writejal(temp, 5'b11111, jalE, writeregE);
	flopenr #(32) hireg3(clk, reset,1, hi, hiE);
	flopenr #(32) loreg3(clk, reset,1, lo, loE);


// Memory stage
	logic [31:0] finalstore;
	flopr #(32) r1M(clk, reset, srcb2E, writedataM);
	flopr #(32) instr2(clk, reset, instrE, instrM);
	flopr #(32) PC2(clk, reset, pcplus4E, pcplus4M);
	flopr #(32) hireg(clk, reset, hiE, hiM);
	flopr #(32) loreg(clk, reset, loE, loM);
	assign sbyte = writedataM[7:0];
	signextbyte seb(sbyte, exsbyte);
	//flopr #(32) ext(clk, reset, exsbyte, exsbyte);
	
//here
	//muxbyte storebyte(tempstore, instrM[1:0], sbyte);
	
	mux2 #(32) WD(writedataM, exsbyte, sbM, finalstore);
	
	flopr #(32) r2M(clk, reset, aluoutE, aluoutM);
	flopr #(5) r3M(clk, reset, writeregE, writeregM);


// Writeback stage
	logic[31:0] finalread;
	flopr #(32) instr3(clk, reset, instrM, instrW);
	flopr #(32) PC3(clk, reset, pcplus4M, pcplus4W);
	flopr #(32) hireg2(clk, reset, hiM, hiW);
	flopr #(32) loreg2(clk, reset, loM, loW);
	flopr #(32) r1W(clk, reset, aluoutM, aluoutW);
	flopr #(32) r2W(clk, reset, readdataM, readdataW);
	flopr #(5) r3W(clk, reset, writeregM, writeregW);
	//muxbyte loadbyte(readdataW, instrW[1:0], lbyte);
	assign lbyte = readdataW[7:0];
	signextbyte leb(lbyte, exlbyte);
	mux2 #(32) RD(readdataW, exlbyte, lbW, finalread);
	
	
	mux4 #(32) resmux(aluoutW, readdataW, loW, hiW, memtoregW,resultW);
	mux2 #(32) wbmux(resultW, pcplus4W, jalregW, resultW);


endmodule



module eqcmp(input logic [31:0] a,b,
	    output logic c);
logic [31:0] x;

	  always @(a or b)
		begin
		c = a==b;
	end
endmodule


module hazard(input logic [4:0] rsD, rtD, rsE, rtE,
		input logic [4:0] writeregE,writeregM, writeregW,
		input logic regwriteE, regwriteM,regwriteW,
		input logic [1:0] memtoregE, memtoregM,
		input logic branchD, bneD,
		output logic forwardaD,forwardbD,
		output logic [1:0] forwardaE, forwardbE,
		output logic stallF, stallD,flushE);

	logic lwstallD, branchstallD;
	
// forwarding sources to D stage (branch equality)
	assign forwardaD = (rsD !=0 & rsD == writeregM &regwriteM);
	assign forwardbD = (rtD !=0 & rtD == writeregM &regwriteM);
// forwarding sources to E stage (ALU)
	always_comb
	begin
	forwardaE = 2'b00; forwardbE = 2'b00;
	if (rsE != 0)
	if (rsE == writeregM & regwriteM)
	forwardaE = 2'b10;
	else if (rsE == writeregW & regwriteW)
	forwardaE = 2'b01;
	if (rtE != 0)
	if (rtE == writeregM & regwriteM)
	forwardbE = 2'b10;
	else if (rtE == writeregW & regwriteW)
	forwardbE = 2'b01;
	end
// stalls
	assign #1 lwstallD = (memtoregE==01) &
	(rtE == rsD | rtE == rtD);
	assign #1 branchstallD = ((branchD | bneD) &(regwriteE &(writeregE == rsD | writeregE == rtD))) | (branchD & ((memtoregM==01) &(writeregM == rsD | writeregM == rtD)));
	assign #1 stallD = lwstallD | branchstallD;
	assign #1 stallF = stallD;
// stalling D stalls all previous stages
	assign #1 flushE = stallD;
// stalling D flushes next stage
// Note: not necessary to stall D stage on store
// if source comes from load;
// instead, another bypass network could
// be added from W to M
endmodule




module floprc #(parameter WIDTH = 8)(input logic clk, reset,clear,
					input logic [WIDTH-1:0] d,
					output logic [WIDTH-1:0] q);
	always_ff @(posedge clk, posedge reset)
		if (reset) q <= #1 0;
	else if (clear) q <= #1 0;
	else q <= #1 d;
endmodule

module flopenrc #(parameter WIDTH = 8)(input logic clk, reset,
					input logic en, clear,
					input logic [WIDTH-1:0] d,
					output logic [WIDTH-1:0] q);
	always_ff @(posedge clk, posedge reset)
		if (reset) q <= #1 0;
		else if (clear) q <= #1 0;
		else if (en) q <= #1 d;
endmodule



module flopr #(parameter WIDTH = 8)
              (input  logic             clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule

module flopenr #(parameter WIDTH = 8)
                (input  logic             clk, reset,
                 input  logic             en,
                 input  logic [WIDTH-1:0] d, 
                 output logic [WIDTH-1:0] q);
 
  always_ff @(posedge clk, posedge reset)
    if      (reset) q <= 0;
    else if (en)    q <= d;
endmodule

module imempipe(input logic [5:0] a,
		output logic [31:0] rd);

	logic [31:0] RAM[63:0];
	initial

	begin
	$readmemh("memfile.dat",RAM);
	end

	assign rd = RAM[a]; // word aligned
endmodule


module dmempipe(input logic clk, we,
	input logic [31:0] a, wd,
	output logic [31:0] rd);
	reg [31:0] RAM[63:0];
	initial
	begin
	$readmemh("memfile.dat",RAM);
	end

	assign rd = RAM[a[31:2]]; // word aligned

	always @(posedge clk)
	if (we)
	RAM[a[31:2]] <= wd;
endmodule



module testbenchpipeall();
	logic clk;
	logic reset;
	logic [31:0] writedata, dataadr;
	logic memwrite;

// instantiate device to be tested
	toppipe dut(clk, reset, writedata, dataadr, memwrite);
// initialize test
	initial
	begin
	reset <= 1; # 10; reset <= 0;
	end
// generate clock to sequence tests
	always
	begin
	clk <= 1; # 5; clk <= 0; # 5;
	end
// check results
	always @(negedge clk)
	begin
	if(memwrite) begin
	if(dataadr === 84 & writedata === 7) begin
	$display("Simulation succeeded");
	$stop;
	end else if (dataadr !== 80) begin
	$display("Simulation failed");
	$stop;
	end
	end
	end
endmodule


module toppipe(input  logic        clk, reset, 
           output logic [31:0] writedata, dataadr, 
           output logic        memwrite);

  	logic [31:0] pc, instr, readdata;
  
  // instantiate processor and memories
  	mipspipe mips(clk, reset, pc, instr, memwrite, dataadr, writedata, readdata);
  	imempipe imem2(pc[7:2], instr);
  	dmempipe dmem(clk, memwrite, dataadr, writedata, readdata);
endmodule




module regfilepipe(input  logic        clk, 
               input  logic        we3, 
               input  logic [4:0]  ra1, ra2, wa3, 
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0];

  // three ported register file
  // read two ports combinationally
  // write third port on rising edge of clk
  // register 0 hardwired to 0
  // note: for pipelined processor, write third port
  // on falling edge of clk

  always_ff @( ~clk)
    if (we3) rf[wa3] <= wd3;	
	
  assign rd1 = (ra1 != 0) ? rf[ra1] : 0;
  assign rd2 = (ra2 != 0) ? rf[ra2] : 0;
endmodule



module ALUpipeall ( a, b, f, shift, y, hi, lo, m);
input logic [31:0] a;
input  logic [31:0] b;
output logic [31:0] y, hi, lo;
input logic [3:0] f;
input logic [4:0] shift;
output logic [63:0] m;

logic [31:0] S, Bout;
 assign Bout = f[2] ? ~b : b;
 assign S = a + Bout + f[2];



/*
000  add
001  sub
010  and
011  or
100  not a
101  xor
110  shift
111  slt
*/
always@(a or b)

case(f)
4'b0000: y <= a & Bout;
4'b0001: y <= a | Bout;
4'b0010: y <= S;
4'b0110: y <= S;
4'b0100: y <= ~a;
4'b0101: y <= (~a&b) | (a&~b);
4'b0110: y <= a - b;
4'b0111: if ((a[31] !== 0) &&  (b[31] !== 1) ) y = 1; else if ((a[31] === b[31] ) && (a[30:0] < b[30:0])) y = 1;  else y = 0;
4'b1000: y <= b << shift;
4'b1001: y <= b >> shift;
4'b1010:
 
	begin
	m = a * b;
	hi = m[63:32]; 
	lo = m[31:0];
	end

4'b1011: 
	begin
	hi <= a % b; 
	lo <= a / b;
	end

endcase

 
endmodule


module alupipe(input logic [31:0] A,input logic[31:0]B,
		   input logic [2:0]alucontrol,
		   output logic [31:0] Y);

 logic [31:0] S, Bout;
 assign Bout = alucontrol[2] ? ~B : B;
 assign S = A + Bout + alucontrol[2];

 always_comb
 case (alucontrol[2:0])
 3'b000: assign Y = A & Bout; //A&B
 3'b001: assign Y = A | Bout; //A|B
 3'b010: assign Y = S; // A + B
 3'b101: assign Y = A | Bout; //A|'B
 3'b110: assign Y = S; // A-B "Gets 2's Complement +1 + A"
 3'b111: assign Y = S[31]; //SLT
 endcase


endmodule

module adder(input  logic [31:0] a, b,
             output logic [31:0] y);

  assign y = a + b;
endmodule

module sl2(input  logic [31:0] a,
           output logic [31:0] y);

  // shift left by 2
  assign y = {a[29:0], 2'b00};
endmodule

module signext(input  logic [15:0] a,
               output logic [31:0] y);
              
  assign y = {{16{a[15]}}, a};
endmodule


module signextbyte( input logic [7:0] a,
			output logic [31:0] b);
	assign b = {{24{a[7]}},a};
endmodule



module flopr #(parameter WIDTH = 8)
              (input  logic             clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule

module flopenr #(parameter WIDTH = 8)
                (input  logic             clk, reset,
                 input  logic             en,
                 input  logic [WIDTH-1:0] d, 
                 output logic [WIDTH-1:0] q);
 
  always_ff @(posedge clk, posedge reset)
    if      (reset) q <= 0;
    else if (en)    q <= d;
endmodule

module mux2 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, 
              input  logic             s, 
              output logic [WIDTH-1:0] y);

  assign y = s ? d1 : d0; 
endmodule

module mux3 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, d2,
              input  logic [1:0]       s, 
              output logic [WIDTH-1:0] y);

  assign #1 y = s[1] ? d2 : (s[0] ? d1 : d0); 
endmodule

module mux4 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, d2, d3,
              input  logic [1:0]       s, 
              output logic [WIDTH-1:0] y);

   always_comb
      case(s)
         2'b00: y <= d0;
         2'b01: y <= d1;
         2'b10: y <= d2;
         2'b11: y <= d3;
      endcase
endmodule

module muxbyte(input  logic [31:0] d,
              input  logic [1:0] s, 
              output logic [7:0] y);

   always_comb
      case(s)
         2'b00: y <= d[7:0];
         2'b01: y <= d[15:8];
         2'b10: y <= d[23:16];
         2'b11: y <= d[31:24];
      endcase
endmodule

